module ALUUNO ( input logic a, b, cin,
                    output logic s, cout);
full_adder full_adder_tres ()
endmodule
